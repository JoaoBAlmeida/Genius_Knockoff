library verilog;
use verilog.vl_types.all;
entity genius_knockoff_vlg_check_tst is
    port(
        arrayed_0_2     : in     vl_logic;
        arrayed_0_1     : in     vl_logic;
        arrayed_0_0     : in     vl_logic;
        arrayed_1_2     : in     vl_logic;
        arrayed_1_1     : in     vl_logic;
        arrayed_1_0     : in     vl_logic;
        arrayed_2_2     : in     vl_logic;
        arrayed_2_1     : in     vl_logic;
        arrayed_2_0     : in     vl_logic;
        arrayed_3_2     : in     vl_logic;
        arrayed_3_1     : in     vl_logic;
        arrayed_3_0     : in     vl_logic;
        arrayed_4_2     : in     vl_logic;
        arrayed_4_1     : in     vl_logic;
        arrayed_4_0     : in     vl_logic;
        arrayed_5_2     : in     vl_logic;
        arrayed_5_1     : in     vl_logic;
        arrayed_5_0     : in     vl_logic;
        arrayed_6_2     : in     vl_logic;
        arrayed_6_1     : in     vl_logic;
        arrayed_6_0     : in     vl_logic;
        arrayed_7_2     : in     vl_logic;
        arrayed_7_1     : in     vl_logic;
        arrayed_7_0     : in     vl_logic;
        arrayed_8_2     : in     vl_logic;
        arrayed_8_1     : in     vl_logic;
        arrayed_8_0     : in     vl_logic;
        arrayed_9_2     : in     vl_logic;
        arrayed_9_1     : in     vl_logic;
        arrayed_9_0     : in     vl_logic;
        arrayed_10_2    : in     vl_logic;
        arrayed_10_1    : in     vl_logic;
        arrayed_10_0    : in     vl_logic;
        arrayed_11_2    : in     vl_logic;
        arrayed_11_1    : in     vl_logic;
        arrayed_11_0    : in     vl_logic;
        arrayed_12_2    : in     vl_logic;
        arrayed_12_1    : in     vl_logic;
        arrayed_12_0    : in     vl_logic;
        arrayed_13_2    : in     vl_logic;
        arrayed_13_1    : in     vl_logic;
        arrayed_13_0    : in     vl_logic;
        arrayed_14_2    : in     vl_logic;
        arrayed_14_1    : in     vl_logic;
        arrayed_14_0    : in     vl_logic;
        arrayed_15_2    : in     vl_logic;
        arrayed_15_1    : in     vl_logic;
        arrayed_15_0    : in     vl_logic;
        arrayed_16_2    : in     vl_logic;
        arrayed_16_1    : in     vl_logic;
        arrayed_16_0    : in     vl_logic;
        arrayed_17_2    : in     vl_logic;
        arrayed_17_1    : in     vl_logic;
        arrayed_17_0    : in     vl_logic;
        arrayed_18_2    : in     vl_logic;
        arrayed_18_1    : in     vl_logic;
        arrayed_18_0    : in     vl_logic;
        arrayed_19_2    : in     vl_logic;
        arrayed_19_1    : in     vl_logic;
        arrayed_19_0    : in     vl_logic;
        arrayed_20_2    : in     vl_logic;
        arrayed_20_1    : in     vl_logic;
        arrayed_20_0    : in     vl_logic;
        arrayed_21_2    : in     vl_logic;
        arrayed_21_1    : in     vl_logic;
        arrayed_21_0    : in     vl_logic;
        arrayed_22_2    : in     vl_logic;
        arrayed_22_1    : in     vl_logic;
        arrayed_22_0    : in     vl_logic;
        arrayed_23_2    : in     vl_logic;
        arrayed_23_1    : in     vl_logic;
        arrayed_23_0    : in     vl_logic;
        arrayed_24_2    : in     vl_logic;
        arrayed_24_1    : in     vl_logic;
        arrayed_24_0    : in     vl_logic;
        led0            : in     vl_logic;
        led1            : in     vl_logic;
        led2            : in     vl_logic;
        led3            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end genius_knockoff_vlg_check_tst;
