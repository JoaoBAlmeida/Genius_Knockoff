library verilog;
use verilog.vl_types.all;
entity genius_knockoff_vlg_vec_tst is
end genius_knockoff_vlg_vec_tst;
