library verilog;
use verilog.vl_types.all;
entity genius_knockoff is
    port(
        clk             : in     vl_logic;
        rst             : in     vl_logic;
        btn0            : in     vl_logic;
        btn1            : in     vl_logic;
        btn2            : in     vl_logic;
        btn3            : in     vl_logic;
        led0            : out    vl_logic;
        led1            : out    vl_logic;
        led2            : out    vl_logic;
        led3            : out    vl_logic;
        arrayed_24_0    : out    vl_logic;
        arrayed_24_1    : out    vl_logic;
        arrayed_24_2    : out    vl_logic;
        arrayed_23_0    : out    vl_logic;
        arrayed_23_1    : out    vl_logic;
        arrayed_23_2    : out    vl_logic;
        arrayed_22_0    : out    vl_logic;
        arrayed_22_1    : out    vl_logic;
        arrayed_22_2    : out    vl_logic;
        arrayed_21_0    : out    vl_logic;
        arrayed_21_1    : out    vl_logic;
        arrayed_21_2    : out    vl_logic;
        arrayed_20_0    : out    vl_logic;
        arrayed_20_1    : out    vl_logic;
        arrayed_20_2    : out    vl_logic;
        arrayed_19_0    : out    vl_logic;
        arrayed_19_1    : out    vl_logic;
        arrayed_19_2    : out    vl_logic;
        arrayed_18_0    : out    vl_logic;
        arrayed_18_1    : out    vl_logic;
        arrayed_18_2    : out    vl_logic;
        arrayed_17_0    : out    vl_logic;
        arrayed_17_1    : out    vl_logic;
        arrayed_17_2    : out    vl_logic;
        arrayed_16_0    : out    vl_logic;
        arrayed_16_1    : out    vl_logic;
        arrayed_16_2    : out    vl_logic;
        arrayed_15_0    : out    vl_logic;
        arrayed_15_1    : out    vl_logic;
        arrayed_15_2    : out    vl_logic;
        arrayed_14_0    : out    vl_logic;
        arrayed_14_1    : out    vl_logic;
        arrayed_14_2    : out    vl_logic;
        arrayed_13_0    : out    vl_logic;
        arrayed_13_1    : out    vl_logic;
        arrayed_13_2    : out    vl_logic;
        arrayed_12_0    : out    vl_logic;
        arrayed_12_1    : out    vl_logic;
        arrayed_12_2    : out    vl_logic;
        arrayed_11_0    : out    vl_logic;
        arrayed_11_1    : out    vl_logic;
        arrayed_11_2    : out    vl_logic;
        arrayed_10_0    : out    vl_logic;
        arrayed_10_1    : out    vl_logic;
        arrayed_10_2    : out    vl_logic;
        arrayed_9_0     : out    vl_logic;
        arrayed_9_1     : out    vl_logic;
        arrayed_9_2     : out    vl_logic;
        arrayed_8_0     : out    vl_logic;
        arrayed_8_1     : out    vl_logic;
        arrayed_8_2     : out    vl_logic;
        arrayed_7_0     : out    vl_logic;
        arrayed_7_1     : out    vl_logic;
        arrayed_7_2     : out    vl_logic;
        arrayed_6_0     : out    vl_logic;
        arrayed_6_1     : out    vl_logic;
        arrayed_6_2     : out    vl_logic;
        arrayed_5_0     : out    vl_logic;
        arrayed_5_1     : out    vl_logic;
        arrayed_5_2     : out    vl_logic;
        arrayed_4_0     : out    vl_logic;
        arrayed_4_1     : out    vl_logic;
        arrayed_4_2     : out    vl_logic;
        arrayed_3_0     : out    vl_logic;
        arrayed_3_1     : out    vl_logic;
        arrayed_3_2     : out    vl_logic;
        arrayed_2_0     : out    vl_logic;
        arrayed_2_1     : out    vl_logic;
        arrayed_2_2     : out    vl_logic;
        arrayed_1_0     : out    vl_logic;
        arrayed_1_1     : out    vl_logic;
        arrayed_1_2     : out    vl_logic;
        arrayed_0_0     : out    vl_logic;
        arrayed_0_1     : out    vl_logic;
        arrayed_0_2     : out    vl_logic
    );
end genius_knockoff;
